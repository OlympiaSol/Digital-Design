library verilog;
use verilog.vl_types.all;
entity REG4_vlg_vec_tst is
end REG4_vlg_vec_tst;
