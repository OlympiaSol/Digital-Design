library verilog;
use verilog.vl_types.all;
entity Reg8Shcematic_vlg_vec_tst is
end Reg8Shcematic_vlg_vec_tst;
