library verilog;
use verilog.vl_types.all;
entity Exercise2_vlg_vec_tst is
end Exercise2_vlg_vec_tst;
