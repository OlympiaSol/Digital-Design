library verilog;
use verilog.vl_types.all;
entity Intro_vlg_vec_tst is
end Intro_vlg_vec_tst;
