library verilog;
use verilog.vl_types.all;
entity Exercise2 is
    port(
        D               : out    vl_logic;
        I3              : in     vl_logic;
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        I1              : in     vl_logic;
        I0              : in     vl_logic;
        I2              : in     vl_logic
    );
end Exercise2;
