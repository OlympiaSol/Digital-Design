library verilog;
use verilog.vl_types.all;
entity Lab1_Exercise1 is
    port(
        Q0              : out    vl_logic;
        PB1             : in     vl_logic;
        PB2             : in     vl_logic;
        Q1              : out    vl_logic;
        Q2              : out    vl_logic;
        Q3              : out    vl_logic
    );
end Lab1_Exercise1;
