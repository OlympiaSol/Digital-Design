library verilog;
use verilog.vl_types.all;
entity Dff_Latchbdf_vlg_vec_tst is
end Dff_Latchbdf_vlg_vec_tst;
