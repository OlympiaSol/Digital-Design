library verilog;
use verilog.vl_types.all;
entity JK_FF_vlg_vec_tst is
end JK_FF_vlg_vec_tst;
