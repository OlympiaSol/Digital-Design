library verilog;
use verilog.vl_types.all;
entity Exercise2_vlg_check_tst is
    port(
        D               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Exercise2_vlg_check_tst;
