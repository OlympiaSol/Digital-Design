library verilog;
use verilog.vl_types.all;
entity MultiplierP_vlg_vec_tst is
end MultiplierP_vlg_vec_tst;
