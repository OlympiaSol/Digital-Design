library verilog;
use verilog.vl_types.all;
entity Exercise3_vlg_vec_tst is
end Exercise3_vlg_vec_tst;
