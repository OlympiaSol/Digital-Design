library verilog;
use verilog.vl_types.all;
entity Exercise3_vlg_sample_tst is
    port(
        I0              : in     vl_logic;
        I1              : in     vl_logic;
        I2              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Exercise3_vlg_sample_tst;
