library verilog;
use verilog.vl_types.all;
entity Exercise4_vlg_vec_tst is
end Exercise4_vlg_vec_tst;
