library verilog;
use verilog.vl_types.all;
entity Counter8Bit_vlg_vec_tst is
end Counter8Bit_vlg_vec_tst;
