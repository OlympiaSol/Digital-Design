library IEEE;
use IEEE.std_logic_1164.all;

entity <entity_name> is
	


	port
	(
		
	);
end <entity_name>;

-- Library Clause(s) (optional)
-- Use Clause(s) (optional)

architecture <arch_name> of <entity_name> is

	-- Declarations (optional)

begin

	-- Process Statement (optional)

	-- Concurrent Procedure Call (optional)

	-- Concurrent Signal Assignment (optional)

	-- Conditional Signal Assignment (optional)

	-- Selected Signal Assignment (optional)

	-- Component Instantiation Statement (optional)

	-- Generate Statement (optional)

end <arch_name>;
