library verilog;
use verilog.vl_types.all;
entity Exercise3_vlg_check_tst is
    port(
        F0              : in     vl_logic;
        F1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Exercise3_vlg_check_tst;
